* XSourceSub. Furnished by dw 23/11/2001.
* subcircuit uses xsource code model
.SUBCKT xsourcesub CLK A1 A2 A3 A4 A5 A6 A7 A8
*

* See DSEQ2 for a sequencer without the built-in clock source.
*Vpulse parameters:   V1   V2   TD   TR   TF  PW  PER 
vclk clk 0 DC 0 pulse (0   5    0    1n   1n  1u  2u)

a1 [Dclk] [D1 D2 D3 D4 D5 D6 D7 D8] dataseq
*
a_dac1 [D1 D2 D3 D4 D5 D6 D7 D8] [A1 A2 A3 A4 A5 A6 A7 A8] dac1
a_adc1 [CLK] [DCLK] adc1
*
.MODEL dataseq xsource(file="{Model_Path}\Misc\XsourceFile.txt" state=[0 5]
+                      strength=[1 1] cycle=40u ttlh=1e-009 tthl=1e-009 vth=1.3)
*
.MODEL dac1 xdac
.MODEL adc1 xadc
*
.ENDS
