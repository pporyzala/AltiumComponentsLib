*Sine of Current
.SUBCKT SINI 1 2 3 4
VX 1 2 0
BX 4 3 I=SIN(I(VX))
.ENDS SINI