*Hyperbolic arc tangent of Current
.SUBCKT ATANHI 1 2 3 4
VX 1 2 0
BX 4 3 I=ATANH(I(VX))
.ENDS ATANHI