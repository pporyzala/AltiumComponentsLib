* Sum relative
* Each input is added to its respective offset and then multiplied by its gain. 
* The results are then summed, multiplied by the output gain and added to the output offset.
* Z = ( ((X2-X1)+offset1)*Gain1 + ((Y2-Y1)+offset2)*Gain2 )* Output Gain + Output Offset
*
* Connections:
*            X1 Positive Input
*            |   X2 Negative Input
*            |   |   Y1 Positive Input
*            |   |   |   Y2 NegativeInput
*            |   |   |   |   Z1 Positive Output
*            |   |   |   |   |   Z2 Negative Output
*            |   |   |   |   |   |
.SUBCKT SUMR 1   2   3   4   5   6 PARAMS: x_offset=0.0 y_offset=0.0 x_gain=1.0 y_gain=1.0 out_gain=1.0 out_offset=0.0
A1 [%vd(1,2) %vd(3,4)] %vd(5,6) sum1
.model sum1 summer(in_offset=[{x_offset} {y_offset}] in_gain=[{x_gain} {y_gain}]
+                  out_gain={out_gain} out_offset={out_offset})
.ENDS SUMR