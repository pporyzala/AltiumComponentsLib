*Hyperbolic arc tangent of Voltage
.SUBCKT ATANHVR 1 2 3 4
BX 3 4 V=ATANH(V(1,2))
.ENDS ATANHVR