*Natural logarithm of Voltage
.SUBCKT LNVR 1 2 3 4
BX 3 4 V=LN(V(1,2))
.ENDS LNVR