*Hyperbolic cosine of Voltage
.SUBCKT COSHV 1 2
BX 2 0 V=COSH(V(1))
.ENDS COSHV