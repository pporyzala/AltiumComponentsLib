*Tangent of Current
.SUBCKT TANI 1 2 3 4
VX 1 2 0
BX 4 3 I=TAN(I(VX))
.ENDS TANI