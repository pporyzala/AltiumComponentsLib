*Square root of Voltage
.SUBCKT SQRTVR 1 2 3 4
BX 3 4 V=SQRT(V(1,2))
.ENDS SQRTVR