*Hyperbolic sine of Current
.SUBCKT SINHI 1 2 3 4
VX 1 2 0
BX 4 3 I=SINH(I(VX))
.ENDS SINHI