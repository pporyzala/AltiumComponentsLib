*Logarithm of Current
.SUBCKT LOGI 1 2 3 4
VX 1 2 0
BX 4 3 I=LOG(I(VX))
.ENDS LOGI