*Natural logarithm of Voltage
.SUBCKT LNV 1 2
BX 2 0 V=LN(V(1))
.ENDS LNV