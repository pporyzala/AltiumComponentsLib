*Arc tangent of Current
.SUBCKT ATANI 1 2 3 4
VX 1 2 0
BX 4 3 I=ATAN(I(VX))
.ENDS ATANI