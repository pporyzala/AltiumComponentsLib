*Hyperbolic arc sine of Current
.SUBCKT ASINHI 1 2 3 4
VX 1 2 0
BX 4 3 I=ASINH(I(VX))
.ENDS ASINHI