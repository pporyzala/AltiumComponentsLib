*Absolute value of Voltage
.SUBCKT ABSV 1 2
BX 2 0 V=ABS(V(1))
.ENDS ABSV