*Hyperbolic arc cosine of Current
.SUBCKT ACOSHI 1 2 3 4
VX 1 2 0
BX 4 3 I=ACOSH(I(VX))
.ENDS ACOSHI