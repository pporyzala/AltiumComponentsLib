* XSourceSub. Furnished by dw 23/11/2001.
* subcircuit uses xsource code model
*
.SUBCKT XSOURCESUB2 A1 A2 A3 A4 A5 A6 A7 A8

A1 [DGND] [D1 D2 D3 D4 D5 D6 D7 D8] DATASEQ

A_ADC1 [0] [DGND] ADC1
A_DAC1 [D1 D2 D3 D4 D5 D6 D7 D8] [A1 A2 A3 A4 A5 A6 A7 A8] DAC1

.MODEL DATASEQ
+ XSOURCE(FILE="D:\Program Files\Design Explorer 99 SE\Library\SIM\MISC\XSOURCEFILE2.TXT" STATE=[0 5] STRENGTH=[1 1] CYCLE=40U TTLH=1E-009 TTHL=1E-009 VTH=1.3)


.MODEL DAC1 XDAC
.MODEL ADC1 XADC

.ENDS