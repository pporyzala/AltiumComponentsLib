*Unary - of Current
.SUBCKT UNARYI 1 2 3 4
VX 1 2 0
BX 4 3 I=-(I(VX))
.ENDS UNARYI