*Sine of Voltage
.SUBCKT SINVR 1 2 3 4
BX 3 4 V=SIN(V(1,2))
.ENDS SINVR