*Exponential of Current
.SUBCKT EXPI 1 2 3 4
VX 1 2 0
BX 4 3 I=EXP(I(VX))
.ENDS EXPI